class Prol16State #(parameter int gRegs = 32);
	pkgProl16::data_v regs[gRegs];
	int programCounter;
	bit cFlag;
	bit zFlag;
	
	function new();
		reset();
	endfunction
	
	task reset();
		for (int i = 0; i < gRegs; i++) begin
			regs[i] = '0;
		end
		programCounter = 0;
		cFlag = 0;
		zFlag = 0;
	endtask
endclass