typedef enum 
	{
		Nop,
		Loadi,
		Jump,
		Jumpc,
		Jumpz,
		Move,
		And,
		Or,
		Xor,
		Not,
		Add,
		Addc,
		Sub,
		Subc,
		Comp,
		Inc,
		Dec,
		Shl,
		Shr,
		Shlc,
		Shrc,
		Invalid
	} Prol16Command;
