package pkgProl16;
	typedef bit [16] data_v;
endpackage