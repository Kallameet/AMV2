class Prol16Opcode;
	int ra;
	int rb;
	Prol16Command cmd;
	data_v data;	
endclass