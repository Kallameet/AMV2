package pkgProl16;
	typedef bit [15:0] data_v;
endpackage
